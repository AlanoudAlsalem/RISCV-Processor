`include "PC.v"
`include "instructionMemory.v"
`include "controlUnit.v"
`include "immGen.v"
`include "registerFile.v"
`include "mux4_1.v"
`include "ALU.v"
`include "dataMemory.v"
`include "mux2_1.v"
`include "branchUnitPred.v"
`include "adder.v"
`include "signExtender.v"
`include "IF_ID.v"
`include "ID_EX.v"
`include "EX_MEM.v"
`include "MEM_WB.v"
`include "forwardingUnit.v"

module microTestbench;
    reg clock;
    reg reset; // reset signal

    // ####################################################### IF #######################################################

    wire PCsrc; // mux selection
    wire [31:0] nextAddress; // mux output

    mux2_1 PCmux(
        .i0(PCplus4),
        .i1(PCjump),
        .select(PCsrc),
        .out(nextAddress)
    );

    wire [31:0] readAddress; // PC output

    PC PC_DUT(
        .nextAddress(nextAddress),
        .clock(clock),
        .reset(reset),
        .nop(nop),
        // when PCsrc = 1 it means that the branch unit is taking the branch
        .branch(PCsrc),
        .readAddress(readAddress)
    );

    wire [31:0] PCplus4, PCjump;

    adder adder1(
        .operand1(readAddress),
        .operand2(32'h4),
        .sum(PCplus4)
    );

    wire [31:0] selectedPCoperand; 

    // supports jalr instruction
    mux2_1 PCadder2(
        .i0(readAddress),
        .i1(ID_forwardedOp1),
        .select(jalr),
        .out(selectedPCoperand)
    );

    adder adder2(
        .operand1(selectedPCoperand),
        .operand2(immediate),
        .sum(PCjump)
    );

    wire [31:0] instruction; // Instruction Memory output
    
    instructionMemory DUT2(
        .instructionAddress(readAddress),
        .instruction(instruction)
    );

    // ####################################################### ID #######################################################

    // IF_ID buffer outputs
    wire [31:0] PC_IF_ID_out, instruction_IF_ID_out;
    wire flush;

    IF_ID buffer1(
        .clock(clock),
        .reset(reset),
        .PC_in(readAddress),
        .instruction_in(instruction),
        .flush(PCsrc),
        // outputs
        .PC(PC_IF_ID_out),
        .instruction(instruction_IF_ID_out)
    );

    wire regWrite, memtoReg, memWrite, sb, lh, ld, jalr, halt; // control signals
    wire [1:0] ALUsrc; // control signal
    wire [3:0] ALUop; // control signal

    controlUnit DUT3(
        .opCode(instruction_IF_ID_out[6:0]),
        .funct3(instruction_IF_ID_out[14:12]),
        .funct7(instruction_IF_ID_out[31:25]),
        .nop(nop),
        .regWrite(regWrite),
        .memtoReg(memtoReg),
        .memWrite(memWrite),
        .ALUsrc(ALUsrc),
        .ALUop(ALUop),
        .sb(sb),
        .lh(lh),
        .ld(ld),
        .jalr(jalr),
        .halt(halt)
    );

    wire [31:0] immediate; // immediate generated by immGen

    immGen DUT4(
        .instruction(instruction_IF_ID_out),
        .out(immediate)
    );

    wire [31:0] readData1, readData2; // Rs1 and Rs2 contents
    wire [31:0] writeData; // WB mux output for reg file
    wire [31:0] r1, r2, r3, r4, r5, r6, r7, r8,
                r9, r10, r11, r12, r13, r14, r15, r16,
                r17, r18, r19, r20, r21, r22, r23, r24,
                r25, r26, r27, r28, r29, r30, r31, r32;

    registerFile DUT5(
        .readReg1(instruction_IF_ID_out[19:15]),
        .readReg2(instruction_IF_ID_out[24:20]),
        .writeReg(rd_MEM_WB_out),
        .writeData(writeData), 
        .regWrite(regWrite_MEM_WB_out),
        .reset(reset),
        .clock(clock),
        .readData1(readData1),
        .readData2(readData2),
        .r1(r1), .r2(r2), .r3(r3), .r4(r4),
        .r5(r5), .r6(r6), .r7(r7), .r8(r8),
        .r9(r9), .r10(r10), .r11(r11), .r12(r12),
        .r13(r13), .r14(r14), .r15(r15), .r16(r16),
        .r17(r17), .r18(r18), .r19(r19), .r20(r20),
        .r21(r21), .r22(r22), .r23(r23), .r24(r24),
        .r25(r25), .r26(r26), .r27(r27), .r28(r28),
        .r29(r29), .r30(r30), .r31(r31), .r32(r32)
    );

    wire [31:0] ID_forwardedOp1, ID_forwardedOp2; // outputs of the two forwarding muxes

    // Rs1 forwarding mux
    mux4_1 fwd1ID(
        .i0(readData1),
        .i1(ALUresult_out), // MEM stage ALU result
        .i2(writeData), // WB stage write result
        .select(ID_forwardOp1),
        .out(ID_forwardedOp1)
    );

    // Rs2 forwarding mux
    mux4_1 fwd2ID(
        .i0(readData2),
        .i1(ALUresult_out), // MEM stage ALU result
        .i2(writeData), // WB stage write result
        .select(ID_forwardOp2),
        .out(ID_forwardedOp2)
    );

    branchUnitPred DUT8(
        .clock(clock),
        .opCode(instruction_IF_ID_out[6:0]),
        .funct3(instruction_IF_ID_out[14:12]),
        .operand1(ID_forwardedOp1),
        .operand2(ID_forwardedOp2),
        .PCsrc(PCsrc)
    );

    // ####################################################### EX #######################################################

    //ID_EX buffer output
    wire regWrite_ID_EX_out, memtoReg_ID_EX_out, sb_ID_EX_out, lh_ID_EX_out;
    wire [1:0] ALUsrc_ID_EX_out;
    wire [3:0] ALUop_ID_EX_out;
    wire [31:0] PC_ID_EX_out, readData1_out, readData2_out, immediate_out;
    wire [4:0] rd_ID_EX_out, rs1, rs2;
    wire ld_ID_EX_out, halt_ID_EX_out;

    ID_EX buffer2(
        .clock(clock),
        .reset(reset),
        .nop(nop),
        // control signals
        .regWrite_in(regWrite),
        .memtoReg_in(memtoReg),
        .memWrite_in(memWrite),
        .sb_in(sb),
        .lh_in(lh),
        .ALUsrc_in(ALUsrc),
        .ALUop_in(ALUop),
        .ld_in(ld),
        .halt_in(halt),
        // PC (address)
        .PC_in(PC_IF_ID_out),
        // registers and immediate
        .readData1_in(readData1),
        .readData2_in(readData2),
        .immediate_in(immediate),
        // register indicies
        .rd_in(instruction_IF_ID_out[11:7]),
        .rs1_in(instruction_IF_ID_out[19:15]),
        .rs2_in(instruction_IF_ID_out[24:20]),

        // outputs
        // control signals
        .regWrite(regWrite_ID_EX_out),
        .memtoReg(memtoReg_ID_EX_out),
        .memWrite(memWrite_ID_EX_out),
        .sb(sb_ID_EX_out),
        .lh(lh_ID_EX_out),
        .ALUsrc(ALUsrc_ID_EX_out),
        .ALUop(ALUop_ID_EX_out),
        .ld(ld_ID_EX_out),
        .halt(halt_ID_EX_out),
        // PC (address)
        .PC(PC_ID_EX_out),
        // registers and immediate
        .readData1(readData1_out),
        .readData2(readData2_out),
        .immediate(immediate_out),
        // register indicies
        .rd(rd_ID_EX_out),
        .rs1(rs1),
        .rs2(rs2)
    );

    wire [1:0] forwardOp1, forwardOp2, ID_forwardOp1, ID_forwardOp2; // MUX selection signals
    wire nop; // nop signal (prevents PC from updating and makes all control signals = 0)

    forwardingUnit DUT1a(
        .clock(clock),
        .reset(reset),
        // opCode from the decode stage (to check for a branch instruction)
        .opCode(instruction_IF_ID_out[6:0]),
        // destination registers from EX MEM and WB stages
        .ID_EX_rd(rd_ID_EX_out),
        .EX_MEM_rd(rd_EX_MEM_out),
        .MEM_WB_rd(rd_MEM_WB_out),
        // source registers from ID and EX stages
        .IF_ID_rs1(instruction_IF_ID_out[19:15]),
        .IF_ID_rs2(instruction_IF_ID_out[24:20]),
        .ID_EX_rs1(rs1),
        .ID_EX_rs2(rs2),
        // regWrite control signal from MEM and WB stage
        .regWrite_EX_MEM(regWrite_EX_MEM_out),
        .regWrite_MEM_WB(regWrite_MEM_WB_out),
        // load signal (load-use hazard)
        .load_ID_EX(ld_ID_EX_out),
        // mux selection signals
        .forwardOp1(forwardOp1),
        .forwardOp2(forwardOp2),
        .ID_forwardOp1(ID_forwardOp1),
        .ID_forwardOp2(ID_forwardOp2),
        // nop for branch and load use hazards
        .nop(nop)
    );

    wire [31:0] rs1Forwarded, rs2Forwarded; // ALU operands after forwarding

    // Rs1 forwarding mux
    mux4_1 fwd1(
        .i0(readData1_out),
        .i1(ALUresult_out), // MEM stage ALU result
        .i2(writeData), // WB stage write result
        .select(forwardOp1),
        .out(rs1Forwarded)
    );

    // Rs2 forwarding mux
    mux4_1 fwd2(
        .i0(readData2_out),
        .i1(ALUresult_out), // MEM stage ALU result
        .i2(writeData), // WB stage write result
        .select(forwardOp2),
        .out(rs2Forwarded)
    );

    wire [31:0] operand2; 

    // choosing the ALU's second operand (register vs immediate vs PC)
    mux4_1 mux2(
        .i0(rs2Forwarded),
        .i1(immediate_out),
        .i2(PC_ID_EX_out),
        .select(ALUsrc_ID_EX_out),
        .out(operand2)
    );

    wire [31:0] ALUresult; // ALU result
    wire zeroFlag; // used in the phase1 version

    ALU DUT6(
        .operation(ALUop_ID_EX_out),
        .operand1(rs1Forwarded),
        .operand2(operand2),
        .result(ALUresult),
        .zeroFlag(zeroFlag)
    );

    // ####################################################### MEM #######################################################

    wire regWrite_EX_MEM_out, memtoReg_out1, memWrite_out1, sb_out1, lh_out1, zeroFlag_out;
    wire [31:0] rs2_out, ALUresult_out;
    wire [4:0] rd_EX_MEM_out;
    wire halt_out1;

    EX_MEM buffer3(
        .clock(clock),
        .reset(reset),
        .regWrite_in(regWrite_ID_EX_out),
        .memtoReg_in(memtoReg_ID_EX_out),
        .memWrite_in(memWrite_ID_EX_out),
        .sb_in(sb_ID_EX_out),
        .lh_in(lh_ID_EX_out),
        .zeroFlag_in(zeroFlag),
        .readData2_in(rs2Forwarded),
        .ALUresult_in(ALUresult),
        .rd_in(rd_ID_EX_out),
        .halt_in(halt_ID_EX_out),
        // outputs
        .regWrite(regWrite_EX_MEM_out),
        .memtoReg(memtoReg_out1),
        .memWrite(memWrite_out1),
        .sb(sb_out1),
        .lh(lh_out1),
        .zeroFlag(zeroFlag_out),
        .readData2(rs2_out),
        .ALUresult(ALUresult_out),
        .rd(rd_EX_MEM_out),
        .halt(halt_out1)
    );

    wire [31:0] data; // data memory output
    wire [31:0] m0,     m4,     m8,     m12,    m16,     
                m20,    m24,    m28,    m32,    m36;

    dataMemory DUT7(
        .dataAddress(ALUresult_out),
        .writeData(rs2_out),
        .memWrite(memWrite_out1),
        .sb(sb_out1),
        .data(data),
        .m0(m0),    .m4(m4),    .m8(m8),    .m12(m12),  .m16(m16),  
        .m20(m20),  .m24(m24),  .m28(m28),  .m32(m32),  .m36(m36)
    );

    wire regWrite_MEM_WB_out, memtoReg_out2, lh_out2;
    wire [31:0] ALUresult_out1, data_out;
    wire [4:0] rd_MEM_WB_out;
    wire halt_out2;

    // ####################################################### WB #######################################################

    MEM_WB buffer4(
        .clock(clock),
        .reset(reset),
        .regWrite_in(regWrite_EX_MEM_out),
        .memtoReg_in(memtoReg_out1),
        .lh_in(lh_out1),
        .ALUresult_in(ALUresult_out),
        .data_in(data),
        .rd_in(rd_EX_MEM_out),
        .halt_in(halt_out1),
        // outputs
        .regWrite(regWrite_MEM_WB_out),
        .memtoReg(memtoReg_out2),
        .lh(lh_out2),
        .ALUresult(ALUresult_out1),
        .data(data_out),
        .rd(rd_MEM_WB_out),
        .halt(halt_out2)
    );

    wire [31:0] outputData;

    signExtender DUT9(
        .lh(lh_out2),
        .inputData(data_out),
        .outputData(outputData)
    );

    mux2_1 mux3(
        .i0(outputData),
        .i1(ALUresult_out1),
        .select(memtoReg_out2),
        .out(writeData)
    );

    // ####################################################### TESTING #######################################################

    initial begin
        clock = 0; reset = 0; #1 reset = 1; #4 reset = 0;
        repeat (20) clock = ~clock;
    end

    integer cycles = 0;

    always @ (posedge clock or posedge halt) begin
        if(halt_out2)
            $finish;
        
        cycles = cycles + 1;
        $display("Cycle #%d", cycles);
        $display("#################### IF ####################");
        $display("selectedPCoperand = %d", selectedPCoperand);
        $display("PC: Next Address = %d Read Address = %d, nop = %b", nextAddress, readAddress, nop);
        $display("IM: Instruction Address= %d Instruction = %h", readAddress, instruction);
        $display("#################### ID ####################");
        $display("CU: opCode = %h, funct3 = %h, funct7 = %h", instruction_IF_ID_out[6:0], instruction_IF_ID_out[14:12], instruction_IF_ID_out[31:25]); 
        $display("nop = %b, regWrite = %b, memtoReg = %b, memWrite = %b, sb = %b, lh = %b, ld = %b, ALUsrc = %b, ALUop = %b, jalr = %b Halt = %b", 
                nop, regWrite, memtoReg, memWrite, sb, lh, ld, ALUsrc, ALUop, jalr, halt);
        $display("IG: immediate = %d", $signed(immediate));
        $display("RF: Rs1 = %d Rs2 = %d", instruction_IF_ID_out[19:15], instruction_IF_ID_out[24:20]);
        $display("Register file content:");
        $display("x0: %d \tx1: %d",   $signed(r1), $signed(r2));
        $display("x2: %d \tx3: %d",   $signed(r3), $signed(r4));
        $display("x4: %d \tx5: %d",   $signed(r5), $signed(r6));
        $display("x6: %d \tx7: %d",   $signed(r7), $signed(r8));
        $display("x8: %d \tx9: %d",   $signed(r9), $signed(r10));
        $display("x10: %d\tx11: %d", $signed(r11), $signed(r12));
        $display("x12: %d\tx13: %d", $signed(r13), $signed(r14));
        $display("x14: %d\tx15: %d", $signed(r15), $signed(r16));
        $display("x16: %d\tx17: %d", $signed(r17), $signed(r18));
        $display("x18: %d\tx19: %d", $signed(r19), $signed(r20));
        $display("x20: %d\tx21: %d", $signed(r21), $signed(r22));
        $display("x22: %d\tx23: %d", $signed(r23), $signed(r24));
        $display("x24: %d\tx25: %d", $signed(r25), $signed(r26));
        $display("x26: %d\tx27: %d", $signed(r27), $signed(r28));
        $display("x28: %d\tx29: %d", $signed(r29), $signed(r30));
        $display("x30: %d\tx31: %d", $signed(r31), $signed(r32));
        $display("ReadData1 = %d ReadData2 = %d", readData1, readData2);
        $display("Branch Unit PCsrc = %b", PCsrc);
        $display("Operand1 = %d, Operand 2 = %d", ID_forwardedOp1, ID_forwardedOp2);
        $display("#################### EX ####################");
        $display("ID_EX_rd = %d EX_MEM_rd = %d MEM_WB_rd = %d", rd_ID_EX_out, rd_EX_MEM_out, rd_MEM_WB_out);
        $display("IF_ID_rs1 = %d IF_ID_rs2 = %d", instruction_IF_ID_out[19:15], instruction_IF_ID_out[24:20]);
        $display("ID_EX_rs1 = %d ID_EX_rs2 = %d", rs1, rs2);
        $display("regWrite EX_MEM = %b regWrite MEM_WB = %b", regWrite_EX_MEM_out, regWrite_MEM_WB_out);
        $display("load = %b", ld_ID_EX_out);
        $display("Forwarding: forwardOp1 = %b forwardOp2 = %b ID_forwardOp1 = %b ID_forwardOp2 = %b nop = %b, opCode = %h", 
            forwardOp1, forwardOp2, ID_forwardOp1, ID_forwardOp2, nop, instruction_IF_ID_out[6:0]);
        $display("ALU: operand 1 = %d operand 2 = %d operation = %h", rs1Forwarded, operand2, ALUop_ID_EX_out);
        $display("Result = %d zeroFlag = %d", ALUresult, zeroFlag);
        $display("#################### MEM ####################");
        $display("Data address = %d, write Data = %d, Data = %d", ALUresult_out, rs2_out, data);
        $display("Data memory contet:");
        $display("m0: %d\tm4: %d", m0, m4);
        $display("m8: %d\tm16: %d", m8, m16);
        $display("m20: %d\tm24: %d", m20, m24);
        $display("m28: %d\tm32: %d", m28, m32);
        $display("m36: %d", m36);
        $display("#################### WB ####################");
        $display("Write data = %d", writeData);
        $display("PCsrc = %b PCplus4 = %d PCjump = %d", PCsrc, PCplus4, PCjump);
        $display("-------------------------------------------------- %t --------------------------------------------------\n", $time);
    end

endmodule
