`include "PC.v"
`include "instructionMemory.v"
`include "controlUnit.v"
`include "immGen.v"
`include "registerFile.v"
`include "mux4_1.v"
`include "ALU.v"
`include "dataMemory.v"
`include "mux2_1.v"
`include "branchUnit.v"
`include "adder.v"

module microTestbench;
    reg clk;
    reg reset; // reset signal

    wire [31:0] nextAddress; // PC input
    wire [31:0] readAddress; // PC output

    wire [31:0] PCplus4, PCjump;

    wire [31:0] instruction; // Instruction Memory output

    wire regWrite, memtoReg, memWrite, sb, halt; // ALU signals
    wire [1:0] ALUsrc; // control signal
    wire [1:0] branch; // control signal
    wire [3:0] ALUop; // control signal

    wire [31:0] immediate; // immediate generated by immGen

    wire [31:0] readData1, readData2; // Rs1 and Rs2

    wire [31:0] operand2; // mux selection

    wire [31:0] ALUresult; // ALU result
    wire zeroFlag;

    wire [31:0] data; // data memory output

    wire [31:0] writeData; // WB mux output for reg file

    wire PCsrc; 

    PC DUT1(
        .nextAddress(nextAddress),
        .clk(clk),
        .reset(reset),
        .readAddress(readAddress)
    );

    adder adder1(
        .operand1(readAddress),
        .operand2(32'h4),
        .sum(PCplus4)
    );

    adder adder2(
        .operand1(readAddress),
        .operand2(immediate),
        .sum(PCjump)
    );

    mux2_1 mux1(
        .i0(PCplus4),
        .i1(PCjump),
        .select(PCsrc),
        .out(nextAddress)
    );
    
    instructionMemory DUT2(
        .instructionAddress(readAddress),
        .instruction(instruction)
    );

    controlUnit DUT3(
        .opCode(instruction[6:0]),
        .funct3(instruction[14:12]),
        .funct7(instruction[31:25]),
        .regWrite(regWrite),
        .memtoReg(memtoReg),
        .memWrite(memWrite),
        .branch(branch),
        .ALUsrc(ALUsrc),
        .ALUop(ALUop),
        .sb(sb),
        .halt(halt)
    );

    immGen DUT4(
        .instruction(instruction),
        .out(immediate)
    );

    registerFile DUT5(
        .readReg1(instruction[19:15]),
        .readReg2(instruction[24:20]),
        .writeReg(instruction[11:7]),
        .writeData(writeData),
        .regWrite(regWrite),
        .reset(reset),
        .readData1(readData1),
        .readData2(readData2)
    );

    mux4_1 mux2(
        .i0(readData1),
        .i1(immediate),
        .i2(readAddress),
        .select(ALUsrc),
        .out(operand2)
    );

    ALU DUT6(
        .operation(ALUop),
        .operand1(readData1),
        .operand2(operand2),
        .result(ALUresult),
        .zeroFlag(zeroFlag)
    );

    dataMemory DUT7(
        .dataAddress(ALUresult),
        .writeData(readData2),
        .memWrite(memWrite),
        .sb(sb),
        .data(data)
    );

    branchUnit DUT8(
        .branch(branch),
        .zeroFlag(zeroFlag),
        .PCsrc(PCsrc)
    );

    mux2_1 mux3(
        .i0(data),
        .i1(ALUresult),
        .select(memtoReg),
        .out(writeData)
    );

    initial begin
        clk = 0; reset = 1; #1 reset = 0; #3
        $display("PC: Next Address = %d Read Address = %d", nextAddress, readAddress);
        $display("IM: Instruction Address= %d Instruction = %h", readAddress, instruction);
        $display("\n");
        $display("CU: opCode = %h, funct7 = %h, funct3 = %h", instruction[6:0], instruction [14:12], instruction [31:25]); 
        $display("regWrite = %b", regWrite);
        $display("memtoReg = %b", memtoReg);
        $display("memWrite = %b", memWrite);
        $display("branch = %b", branch);
        $display("sb = %b", sb);
        $display("ALUsrc = %b", ALUsrc);
        $display("ALUop = %b", ALUop);
        $display("Halt = %b", halt);
        $display("\n");
        $display("IG: immediate = %d", immediate);
        $display("RF: Rs1 = %d Rs2 = %d", readData1, readData2);
        $display("ALU: operand 1 = %d operand 2 = %d operation = %h", readData1, operand2, ALUop);
        $display("Result = %d zeroFlag = %d", ALUresult, zeroFlag);
        $display("Data address = %d, write Data = %d", ALUresult, readData2);
        $display("Data = %d", data);
        $display("\n");
        $display("Write data = %d", writeData);
        $display("PCsrc = %b", PCsrc);
        $display("PCplus4 = %d PCjump = %d", PCplus4, PCjump);

        $display(" %t ------------------------------\n", $time);

        clk = ~clk; #3

        $display("PC: Next Address = %d Read Address = %d", nextAddress, readAddress);
        $display("IM: Instruction Address= %d Instruction = %h", readAddress, instruction);
        $display("\n");
        $display("CU: opCode = %h, funct7 = %h, funct3 = %h", instruction[6:0], instruction [14:12], instruction [31:25]); 
        $display("regWrite = %b", regWrite);
        $display("memtoReg = %b", memtoReg);
        $display("memWrite = %b", memWrite);
        $display("branch = %b", branch);
        $display("sb = %b", sb);
        $display("ALUsrc = %b", ALUsrc);
        $display("ALUop = %b", ALUop);
        $display("Halt = %b", halt);
        $display("\n");
        $display("IG: immediate = %d", immediate);
        $display("RF: Rs1 = %d Rs2 = %d", readData1, readData2);
        $display("ALU: operand 1 = %d operand 2 = %d operation = %h", readData1, operand2, ALUop);
        $display("Result = %d zeroFlag = %d", ALUresult, zeroFlag);
        $display("Data address = %d, write Data = %d", ALUresult, readData2);
        $display("Data = %d", data);
        $display("\n");
        $display("Write data = %d", writeData);
        $display("Write reg = %d", instruction[11:7]);
        $display("PCsrc = %b", PCsrc);
        $display("PCplus4 = %d PCjump = %d", PCplus4, PCjump);
        
        $display(" %t ------------------------------\n", $time);
        clk = ~clk; #1
        clk = ~clk; #3
        $display("PC: Next Address = %d Read Address = %d", nextAddress, readAddress);
        $display("IM: Instruction Address= %d Instruction = %h", readAddress, instruction);
        $display("\n");
        $display("CU: opCode = %h, funct7 = %h, funct3 = %h", instruction[6:0], instruction [14:12], instruction [31:25]); 
        $display("regWrite = %b", regWrite);
        $display("memtoReg = %b", memtoReg);
        $display("memWrite = %b", memWrite);
        $display("branch = %b", branch);
        $display("sb = %b", sb);
        $display("ALUsrc = %b", ALUsrc);
        $display("ALUop = %b", ALUop);
        $display("Halt = %b", halt);
        $display("\n");
        $display("IG: immediate = %d", immediate);
        $display("RF: Rs1 = %d Rs2 = %d", readData1, readData2);
        $display("ALU: operand 1 = %d operand 2 = %d operation = %h", readData1, operand2, ALUop);
        $display("Result = %d zeroFlag = %d", ALUresult, zeroFlag);
        $display("Data address = %d, write Data = %d", ALUresult, readData2);
        $display("Data = %d", data);
        $display("\n");
        $display("Write data = %d", writeData);
        $display("Write reg = %d", instruction[11:7]);
        $display("PCsrc = %b", PCsrc);
        $display("PCplus4 = %d PCjump = %d", PCplus4, PCjump);
        
        $display(" %t ------------------------------\n", $time);
    end

endmodule
