// The interconnection of all components to form the CPU

module CPU(

);

endmodule